module MMIO(
    input clk,
    input wire [11:0] addr,
    input wire mwe,
    input wire [31:0] data,
    output wire [31:0] data_out,
    input wire BTNU,
    output reg  [3:0]  texture_idx
);
    always @(posedge clk) begin
        if (mwe) begin
            case (addr)
                12'd1001: texture_idx <= data[3:0]; 
            endcase
        end
    end

    assign data_out = (addr == 1000) ? {31'b0, BTNU} :
                    (addr == 1001) ? {28'b0, texture_idx} :
                    data;
endmodule
