module and_32 (A, B, Y);
	input  [31:0] A;
	input  [31:0] B;
	output [31:0] Y;

	genvar i;
	generate
		for (i = 0; i<32; i = i + 1) begin: and32
			and (Y[i], A[i], B[i]);
		end
	endgenerate
endmodule

